module test(
	input clk,
	output clk_div
	);
	reg [3:0] count=0;
endmodule

