module test(
	input clk,
	output clk_div
	);
endmodule
